module Color_Palette (
    input [3:0] index,
    output [11:0] RGB_Color
);

    always_comb begin
        // replace with case statement:
      
    end
endmodule